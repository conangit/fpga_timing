
module pipeline_booth_multiplier(
    clk,
    a,
    b,
    product
    );
    
    input clk;
    input [7:0]a;
    input [7:0]b;
    output [15:0]product;
    
    /***************************/
    
    reg [16:0]p[8:0]; //booth算法需要9个步骤
    reg [15:0]item[7:0]; //每个计算步骤(共8个)都有固定的a和a的取反加1
    reg [7:0]diff1[7:0];
    reg [7:0]diff2[7:0];
    
    always @(posedge clk) begin
        /***************************/ //init step
        p[0] <= {8'd0, b, 1'b0};
        item[0] <= {~a + 1'b1, a};
        
        /***************************/ //step 0
        diff1[0] = p[0][16:9] + item[0][7:0];
        diff2[0] = p[0][16:9] + item[0][15:8];
        
        if (p[0][1:0] == 2'b01)
            p[1] <= {diff1[0][7], diff1[0], p[0][8:1]};
        else if (p[0][1:0] == 2'b10)
            p[1] <= {diff2[0][7], diff2[0], p[0][8:1]};
        else
            p[1] <= {p[0][16], p[0][16:1]};
            
        item[1] <= item[0];
        
        /***************************/ //step 1
        diff1[1] = p[1][16:9] + item[1][7:0];
        diff2[1] = p[1][16:9] + item[1][15:8];
        
        if (p[1][1:0] == 2'b01)
            p[2] <= {diff1[1][7], diff1[1], p[1][8:1]};
        else if (p[1][1:0] == 2'b10)
            p[2] <= {diff2[1][7], diff2[1], p[1][8:1]};
        else
            p[2] <= {p[1][16], p[1][16:1]};
            
        item[2] <= item[1];
        
        /***************************/ //step 2
        diff1[2] = p[2][16:9] + item[2][7:0];
        diff2[2] = p[2][16:9] + item[2][15:8];
        
        if (p[2][1:0] == 2'b01)
            p[3] <= {diff1[2][7], diff1[2], p[2][8:1]};
        else if (p[2][1:0] == 2'b10)
            p[3] <= {diff2[2][7], diff2[2], p[2][8:1]};
        else
            p[3] <= {p[2][16], p[2][16:1]};
            
        item[3] <= item[2];
        
        /***************************/ //step 3
        diff1[3] = p[3][16:9] + item[3][7:0];
        diff2[3] = p[3][16:9] + item[3][15:8];
        
        if (p[3][1:0] == 2'b01)
            p[4] <= {diff1[3][7], diff1[3], p[3][8:1]};
        else if (p[3][1:0] == 2'b10)
            p[4] <= {diff2[3][7], diff2[3], p[3][8:1]};
        else
            p[4] <= {p[3][16], p[3][16:1]};
            
        item[4] <= item[3];
       
        /***************************/ //step 4
        diff1[4] = p[4][16:9] + item[4][7:0];
        diff2[4] = p[4][16:9] + item[4][15:8];
        
        if (p[4][1:0] == 2'b01)
            p[5] <= {diff1[4][7], diff1[4], p[4][8:1]};
        else if (p[4][1:0] == 2'b10)
            p[5] <= {diff2[4][7], diff2[4], p[4][8:1]};
        else
            p[5] <= {p[4][16], p[4][16:1]};
            
        item[5] <= item[4];
       
        /***************************/ //step 5
        diff1[5] = p[5][16:9] + item[5][7:0];
        diff2[5] = p[5][16:9] + item[5][15:8];
        
        if (p[5][1:0] == 2'b01)
            p[6] <= {diff1[5][7], diff1[5], p[5][8:1]};
        else if (p[5][1:0] == 2'b10)
            p[6] <= {diff2[5][7], diff2[5], p[5][8:1]};
        else
            p[6] <= {p[5][16], p[5][16:1]};
            
        item[6] <= item[5];
        
        /***************************/ //step 6
        diff1[6] = p[6][16:9] + item[6][7:0];
        diff2[6] = p[6][16:9] + item[6][15:8];
        
        if (p[6][1:0] == 2'b01)
            p[7] <= {diff1[6][7], diff1[6], p[6][8:1]};
        else if (p[6][1:0] == 2'b10)
            p[7] <= {diff2[6][7], diff2[6], p[6][8:1]};
        else
            p[7] <= {p[6][16], p[6][16:1]};
            
        item[7] <= item[6];
        
        /***************************/ //step 7
        diff1[7] = p[7][16:9] + item[7][7:0];
        diff2[7] = p[7][16:9] + item[7][15:8];
        
        if (p[7][1:0] == 2'b01)
            p[8] <= {diff1[7][7], diff1[7], p[7][8:1]};
        else if (p[7][1:0] == 2'b10)
            p[8] <= {diff2[7][7], diff2[7], p[7][8:1]};
        else
            p[8] <= {p[7][16], p[7][16:1]};
            
        // item[8] <= item[7];
    end
    
    assign product = p[8][16:1];
    
    
endmodule


